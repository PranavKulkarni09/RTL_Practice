module model #(parameter
  DATA_WIDTH = 16
) (
  input [DATA_WIDTH-1:0] din,
  output logic [$clog2(DATA_WIDTH):0] dout
);

  logic [$clog2(DATA_WIDTH):0] temp;

  always @ (*) begin
    temp = 0;
    for(int i = 0; i<DATA_WIDTH; i++) begin
      if(din[i]==1)begin
        temp++;
      end
    end
    dout = temp;
  end

endmodule
